***** Spice Netlist for Cell 'invX1' *****

************** Module invX1 **************
.subckt invX1 in out
m0 out in gnd gnd scmosn w='0.6u' l='0.4u' m='1' 
m1 out in vdd vdd scmosp w='0.6u' l='0.4u' m='1' 
.ends invX1


.end

